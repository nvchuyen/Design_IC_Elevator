module scan_kbcode
	( 	
		input wire clk , reset, 
		input wire ps2d, ps2c, rd_en,
		output wire [7:0] key_code  
	);

	localparam BRK = 8'hf0; // break code 
// symbolic state declaration 
	localparam 	wait_brk = 1'b0, 
					get_code = 1'b1;
					
// signal declaration 
	reg state_reg , state_next; 
	wire [7:0] scan_out ; 
	wire scan_done_tick;
	reg got;	
	
	ps2_rx ps2_unit 
	(
		.clk (clk), 
		.reset (reset), 
		.rx_en (1'b1), 																						
		.ps2d (ps2d), 
		.ps2c (ps2c), 
		.rx_done_tick (scan_done_tick), 
		.dout (scan_out)
	);
	
	memory r1
	(
		.clk (clk),
		.reset(reset),	
		.wr_en (got), 
		.data_in (scan_out),
		.q(key_code)
	);
	always @(posedge clk, posedge reset) 
		if (reset ) 
			state_reg <= wait_brk ; 
		else
			if(~rd_en)
				state_reg <= wait_brk ;
			else	
				state_reg <= state_next ; 

	always@(*) 
	begin
		got = 1'b0;
		state_next = state_reg; 
		
		case (state_reg) 
			wait_brk: // wait for FO of break code 
				if (scan_done_tick == 1'b1 && scan_out == BRK) 
					state_next = get_code ;
					
			get_code: // get the following scan code 
				if (scan_done_tick) 
				begin 
					got = 1'b1; 
					state_next = wait_brk ; 
				end
		endcase	
	end
endmodule
